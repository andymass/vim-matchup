module somemodule
always@( * ) begin
    //begin
end

///end
endmodule
